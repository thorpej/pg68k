/*
 * Copyright (c) 2025 Jason R. Thorpe.
 * All rights reserved.
 *
 * Redistribution and use in source and binary forms, with or without
 * modification, are permitted provided that the following conditions
 * are met:
 * 1. Redistributions of source code must retain the above copyright
 *    notice, this list of conditions and the following disclaimer.
 * 2. Redistributions in binary form must reproduce the above copyright
 *    notice, this list of conditions and the following disclaimer in the
 *    documentation and/or other materials provided with the distribution.
 *
 * THIS SOFTWARE IS PROVIDED BY THE AUTHOR ``AS IS'' AND ANY EXPRESS OR
 * IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES
 * OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.
 * IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR ANY DIRECT, INDIRECT,
 * INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING,
 * BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
 * LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED
 * AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
 * OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
 * OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
 * SUCH DAMAGE.
 */

/*
 * Playground 68030 System Controller.
 *
 * This contains most of the random glue logic, top-level address
 * decoding, fast-RAM memory interface, and bus error generation.
 */

module sysctl(
	input wire nRST,
	input wire DRAM_CLK,

	input wire nAS,
	input wire nDS,
	input wire RnW,
	input wire [1:0] SIZ,

	input wire [2:0] FC,
	input wire [31:0] ADDR,

	input wire nCBREQ,

	output wire STERM,		/* external open-drain inv */
	output wire CI,			/* external open-drain inv */
	output wire CBACK,		/* external open-drain inv */
	output wire BERR,		/* external open-drain inv */
	output wire [1:0] DSACK,	/* external open-drain inv */

	output wire nROMSEL,
	output wire nEXPSEL,
	output wire [3:0] nDRAMSEL,
	output wire nFPUSEL,
	output wire nIACKSEL,

	output wire nISASEL,
	output wire nPSUCSEL,
	output wire nINTCSEL,
	output wire nI2CSEL,

	output wire CPU_CLK,
	output wire CLK_6_25,

	output wire nFRAMSEL,
	output wire nFRAM_RD,
	output wire nFRAM_WR,
	output wire [3:0] nFRAM_BE,

	output wire RESET
);

/*
 * Clock generation.  We receive the DRAM clock as input (50MHz).  We
 * produce the following clock outputs:
 *
 * - CPU_CLK (25MHz)	DRAM_CLK / 2
 * - CLK_6_25 (6.25MHz)	DRAM_CLK / 8
 */
reg [2:0] ClockDivider;
always @(posedge DRAM_CLK) begin
//
// We want the clock to be already free-running and stable when other
// devices come out of reset, so do not reset the counter.  The power-
// on-reset is elongated to ensure many cycles of free-running before
// other devices begin consuming it.
//
//	if (~nRST)
//		ClockDivider <= 3'd0;
//	else
		ClockDivider <= ClockDivider + 3'd1;
end
assign CPU_CLK = ClockDivider[0];
assign CLK_6_25 = ClockDivider[2];

/*
 * We count the first 4 bus cycles after a /RESET occurs, and use that
 * to ensure the ROM is selected for the reset vector fetch.
 *
 * N.B. We want the state to advance **after** the bus cycle is over,
 * thus we clock on the rising edge of nAS.
 */
reg [1:0] BootState;
always @(posedge nAS, negedge nRST) begin
	if (~nRST)
		BootState <= 2'd0;
	else begin
		if (BootState != 2'd3)
			BootState <= BootState + 2'd1;
	end
end
wire ResetVecFetch;
assign ResetVecFetch = (BootState != 2'd3);

/*
 * Bus error generation.
 *
 * This will drive the BERR output to the CPU if a bus cycle fails
 * to terminate after 64 CPU clock cycles.
 *
 * If /RESET is asserted or there is not active bus cycle (/AS not asserted),
 * then we reset the counter to 0.
 *
 * No other termination indication is required other than de-assertion of
 * /AS; when bus cycles terminate by whatever means, the CPU de-asserts /AS
 * before the rising edge of the CPU clock cycle that begins the next bus
 * cycle's S0.
 */
reg [5:0] BerrState;
always @(posedge CPU_CLK, negedge nRST) begin
	if (~nRST)
		BerrState <= 6'd0;
	else begin
		if (nAS)
			BerrState <= 6'd0;
		else if (BerrState != 6'd63)
			BerrState <= BerrState + 6'd1;
	end
end
assign BERR = (BerrState == 6'd63);

/*
 * Function bits for address space encodings:
 *
 * FC2   FC1   FC0
 *  0     0     0       (Undefined, reserved)
 *  0     0     1       User Data Space
 *  0     1     0       User Program Space
 *  0     1     1       (Undefined, reserved)
 *  1     0     0       (Undefined, reserved)
 *  1     0     1       Supervisor Data Space
 *  1     1     0       Supervisor Program Space
 *  1     1     1       CPU Space
 *
 * Note that {User,Supervisor}{Data,Program} -> FC1 xor FC0 -> 1
 */
wire SpaceNormal = (FC[1] ^ FC[0]);
wire SpaceCPU = (FC == 3'd7);

localparam QUAL_nAS	= 2'bx0;
localparam QUAL_nCLK	= 2'b0x;
wire [1:0] AddrQual = {CPU_CLK, nAS};

localparam SPC_CPU	= 2'b10;
localparam SPC_NORM	= 2'b01;
wire [1:0] AddrSpace = {SpaceCPU, SpaceNormal};

/*
 * Top-level address decoding:
 *
 * $FFF0.0000 - $FFFF.FFFF      System ROM (1MB)
 * $FFE0.0000 - $FFEF.FFFF      Peripheral device space (1MB)
 *     0.0000 -     0.FFFF	  (ISA I/O space)
 * $FE00.0000 - $FE3F.FFFF      Fast RAM (4MB)
 * $8000.0000 - $80FF.FFFF      Expansion space (16MB)
 * $0000.0000 - $3FFF.FFFF      DRAM (1GB, as 4x256MB)
 *
 * The DRAM region is arranged as up-to-four discrete 256MB banks, each
 * controlled by a DRAMCTL.
 *
 * Expansion space is further decoded externally, qualified by /EXPSEL.
 *
 * The peripheral space is divided into two regions, one with ISA-like
 * peripherals externally decoded and qualified by /ISASEL, and other
 * on-board peripherals that speak the native 68030 bus protocol decoded
 * below.
 */

/*			          Address bits
 *			      31               13
 *			      |                 |			*/
localparam REGION_ROM	= 19'b111111111111xxxxxxx;
localparam REGION_DEV	= 19'b111111111110xxxxxxx;
/*         REGION_FRAM	= 19'b1111111000xxxxxxxxx; Handled below.	*/
localparam REGION_EXP	= 19'b10000000xxxxxxxxxxx;
localparam REGION_DRAM0	= 19'b0000xxxxxxxxxxxxxxx;
localparam REGION_DRAM1	= 19'b0001xxxxxxxxxxxxxxx;
localparam REGION_DRAM2	= 19'b0010xxxxxxxxxxxxxxx;
localparam REGION_DRAM3	= 19'b0011xxxxxxxxxxxxxxx;

	/* (CPU space) ACCTYPE = 0x02 (coproc), CPID = 0x01 */
localparam REGION_FPU	= 19'bxxxxxxxxxxxx0010001;

	/* (CPU space) ACCTYPE = 0x0f (IACK) */
localparam REGION_IACK	= 19'bxxxxxxxxxxxx1111xxx;

localparam RV_Y		= 1'b1;
localparam RV_N		= 1'b0;
localparam RV_X		= 1'bx;

localparam SEL_NONE	= 9'b111111111;
localparam SEL_ROM	= 9'b111111110;
localparam SEL_DEV	= 9'b111111101;
localparam SEL_EXP	= 9'b111111011;
localparam SEL_DRAM0	= 9'b111110111;
localparam SEL_DRAM1	= 9'b111101111;
localparam SEL_DRAM2	= 9'b111011111;
localparam SEL_DRAM3	= 9'b110111111;
localparam SEL_FPU	= 9'b101111111;
localparam SEL_IACK	= 9'b011111111;

wire nDEVSELx;
wire nROMSELx;
reg [8:0] SelectOutputs;
always @(*) begin
	casex ({AddrQual, AddrSpace, ResetVecFetch, ADDR[31:13]})
	{QUAL_nAS,  SPC_NORM, RV_X, REGION_ROM}:   SelectOutputs = SEL_ROM;

	{QUAL_nAS,  SPC_NORM, RV_X, REGION_DEV}:   SelectOutputs = SEL_DEV;

	{QUAL_nAS,  SPC_NORM, RV_X, REGION_EXP}:   SelectOutputs = SEL_EXP;

	{QUAL_nAS,  SPC_NORM, RV_Y, REGION_DRAM0}: SelectOutputs = SEL_ROM;
	{QUAL_nAS,  SPC_NORM, RV_N, REGION_DRAM0}: SelectOutputs = SEL_DRAM0;
	{QUAL_nAS,  SPC_NORM, RV_X, REGION_DRAM1}: SelectOutputs = SEL_DRAM1;
	{QUAL_nAS,  SPC_NORM, RV_X, REGION_DRAM2}: SelectOutputs = SEL_DRAM2;
	{QUAL_nAS,  SPC_NORM, RV_X, REGION_DRAM3}: SelectOutputs = SEL_DRAM3;

	{QUAL_nCLK, SPC_CPU,  RV_X, REGION_FPU}:   SelectOutputs = SEL_FPU;
	{QUAL_nAS,  SPC_CPU,  RV_X, REGION_FPU}:   SelectOutputs = SEL_FPU;

	{QUAL_nAS,  SPC_CPU,  RV_X, REGION_IACK}:  SelectOutputs = SEL_IACK;

	default:                                   SelectOutputs = SEL_NONE;
	endcase
end
assign {nIACKSEL, nFPUSEL, nDRAMSEL, nEXPSEL, nDEVSELx, nROMSELx}
    = SelectOutputs;

/*
 * ROM only selected for read cycles.  /ROMSEL can be connected to /CS
 * and /OE on both of the SST39SF040-70s.
 */
assign nROMSEL = nROMSELx | ~RnW;

/*
 * Further qualify the DEV space:
 *
 * 0.xxxx	ISA I/O space
 *			(DUART, Timer, ATA disk, Ethernet)
 * 1.000x	PCF8584 I2C controller
 * F.FFEx	PSU controller
 * F.FFFx	Interrupt controller
 */
localparam DEV_ISA	= 20'h0xxxx;
localparam DEV_I2C	= 20'h1000x;
localparam DEV_PSUC	= 20'hFFFEx;
localparam DEV_INTC	= 20'hFFFFx;

localparam DSEL_NONE	= 4'b1111;
localparam DSEL_ISA	= 4'b0111;
localparam DSEL_I2C	= 4'b1011;
localparam DSEL_PSUC	= 4'b1101;
localparam DSEL_INTC	= 4'b1110;

reg [2:0] DevSelectOutputs;
always @(*) begin
	casex ({nDEVSELx, nDS, RnW, ADDR[19:0]})
	{1'b0, 1'bx, 1'bx, DEV_ISA}:  DevSelectOutputs = DSEL_ISA;
	/*
	 * The PSU controller is wired up so that any time it is
	 * selected, it will either reset or power off the system
	 * (depending on the value of D0).  So, avoid errant reads,
	 * and only select it once the data bus is valid.
	 */
	{1'b0, 1'b0, 1'b0, DEV_PSUC}: DevSelectOutputs = DSEL_PSUC;
	{1'b0, 1'bx, 1'bx, DEV_INTC}: DevSelectOutputs = DSEL_INTC;
	/*
	 * Also need to qual /I2CSEL on /DS because we want to
	 * ensure that the PCF8584 comes up in 68000 interface
	 * mode.
	 */
	{1'b0, 1'b0, 1'bx, DEV_I2C}:  DevSelectOutputs = DSEL_I2C;
	default:                      DevSelectOutputs = DSEL_NONE;
	endcase
end
assign {nISASEL, nI2CSEL, nPSUCSEL, nINTCSEL}
    = DevSelectOutputs;

localparam REGION_FRAM = 10'b1111111100;

/* 
 *           nFRAM_BE[3:0] ------++
 *                nFRAM_WR ----+ ||
 *                nFRAM_RD ---+| ||
 *                   STERM --+|| ||
 *                           |||-++-				*/
localparam FRS_NONE	= 7'b0111111;

localparam FRS_RD	= 7'b1011111;

localparam FRS_WR1_0	= 7'b1100111;
localparam FRS_WR1_1	= 7'b1101011;
localparam FRS_WR1_2	= 7'b1101101;
localparam FRS_WR1_3	= 7'b1101110;

localparam FRS_WR2_0	= 7'b1100011;
localparam FRS_WR2_1	= 7'b1101001;
localparam FRS_WR2_2	= 7'b1101100;
localparam FRS_WR2_3	= 7'b1101110;

localparam FRS_WR3_0	= 7'b1100001;
localparam FRS_WR3_1	= 7'b1101000;
localparam FRS_WR3_2	= 7'b1101100;
localparam FRS_WR3_3	= 7'b1101110;

localparam FRS_WR4_0	= 7'b1100000;
localparam FRS_WR4_1	= 7'b1101000;
localparam FRS_WR4_2	= 7'b1101100;
localparam FRS_WR4_3	= 7'b1101110;

reg [6:0] FRSOutputs;
always @(*) begin
	casex ({nAS, AddrSpace, ADDR[31:22], RnW, SIZ[1:0], ADDR[1:0]})
	/*
	 * Byte enables, from Table 7-4 in the 68030 User's Manual.
	 * N.B. for reads, we enable all bytes.
	 */

	/* reads */
	{1'b0, SPC_NORM, REGION_FRAM, 5'b1xxxx}:  FRSOutputs = FRS_RD;

	/* byte writes */
	{1'b0, SPC_NORM, REGION_FRAM, 5'b00100}:  FRSOutputs = FRS_WR1_0;
	{1'b0, SPC_NORM, REGION_FRAM, 5'b00101}:  FRSOutputs = FRS_WR1_1;
	{1'b0, SPC_NORM, REGION_FRAM, 5'b00110}:  FRSOutputs = FRS_WR1_2;
	{1'b0, SPC_NORM, REGION_FRAM, 5'b00111}:  FRSOutputs = FRS_WR1_3;

	/* word writes */
	{1'b0, SPC_NORM, REGION_FRAM, 5'b01000}:  FRSOutputs = FRS_WR2_0;
	{1'b0, SPC_NORM, REGION_FRAM, 5'b01001}:  FRSOutputs = FRS_WR2_1;
	{1'b0, SPC_NORM, REGION_FRAM, 5'b01010}:  FRSOutputs = FRS_WR2_2;
	{1'b0, SPC_NORM, REGION_FRAM, 5'b01011}:  FRSOutputs = FRS_WR2_3;

	/* 3 byte writes */
	{1'b0, SPC_NORM, REGION_FRAM, 5'b01100}:  FRSOutputs = FRS_WR3_0;
	{1'b0, SPC_NORM, REGION_FRAM, 5'b01101}:  FRSOutputs = FRS_WR3_1;
	{1'b0, SPC_NORM, REGION_FRAM, 5'b01110}:  FRSOutputs = FRS_WR3_2;
	{1'b0, SPC_NORM, REGION_FRAM, 5'b01111}:  FRSOutputs = FRS_WR3_3;

	/* long word writes */
	{1'b0, SPC_NORM, REGION_FRAM, 5'b00000}:  FRSOutputs = FRS_WR4_0;
	{1'b0, SPC_NORM, REGION_FRAM, 5'b00001}:  FRSOutputs = FRS_WR4_1;
	{1'b0, SPC_NORM, REGION_FRAM, 5'b00010}:  FRSOutputs = FRS_WR4_2;
	{1'b0, SPC_NORM, REGION_FRAM, 5'b00011}:  FRSOutputs = FRS_WR4_3;

	default:                                  FRSOutputs = FRS_NONE;
	endcase
end
assign {STERM, nFRAM_RD, nFRAM_WR, nFRAM_BE} = FRSOutputs;
assign nFRAMSEL = ~STERM;	/* we only assert STERM for Fast RAM */
assign CBACK = 1'b0;

/* Inhibit cache if fetching the reset vector or accessing DEV space. */
assign CI = (ResetVecFetch || ~nDEVSELx);

/*
 * Bus cycle state machine.
 *
 * Generate DSACKx based on the selected device and its timing constraints.
 *
 * Note we only do this for devices that don't do the 68000 bus protocol
 * natively, which means: the ROM.  (ISA devices are handled by the ISA
 * controller.)
 */
reg [1:0] dsack;
localparam PORT_1	= 2'b01;
localparam PORT_2	= 2'b10;

reg [1:0] BCState;
localparam BC_Idle	= 4'd0;
localparam BC_B1W1	= 4'd1;	/* bytes: 1, waits: 1 */
localparam BC_B2W1	= 4'd2;	/* bytes: 2, waits: 1 */
localparam BC_Finish	= 4'd3;

always @(posedge CPU_CLK, negedge nRST) begin
	if (~nRST) begin
		BCState <= 2'd0;
		dsack <= 2'b00;
	end
	else begin
		case (BCState)
		BC_Idle: begin
			if (~nROMSEL) begin
				/*
				 * /ROMSEL is doing all the work required,
				 * but we need 1 wait state to meet the
				 * 70ns access time.
				 */
				BCState <= BC_B2W1;
			end
			else if (~nPSUCSEL) begin
				/*
				 * Writing to the PSU controller will
				 * either reset or power off the system,
				 * and it does not participate in the
				 * bus protocol whatsoever.  Just provide
				 * a single wait-state to make sure D0 is
				 * stable in the latch fronting the
				 * microcontroller, and then terminate
				 * the bus cycle.  The system will reset
				 * or power off a few milliseconds later.
				 */
				BCState <= BC_B1W1;
			end
		end

		BC_B1W1: begin
			dsack <= PORT_1;
			BCState <= BC_Finish;
		end

		BC_B2W1: begin
			dsack <= PORT_2;
			BCState <= BC_Finish;
		end

		BC_Finish: begin
			if (nDS) begin
				dsack <= 2'b00;
				BCState <= BC_Idle;
			end
		end
		endcase
	end
end

/*
 * Qual with /DS from the CPU so they de-assert immediately.
 */
assign DSACK = dsack & {~nDS, ~nDS};

/* Generate a positive-level reset signal for anything that needs it. */
assign RESET = ~nRST;

endmodule

// Pin assignment for Yosys workflow.
//
//PIN: CHIP "sysctl" ASSIGNED TO AN TQFP100
//
//     === Inputs ===
//PIN: nCBREQ		: 30
//PIN: RnW		: 31
//PIN: SIZ_0		: 32
//PIN: SIZ_1		: 33
//PIN: ADDR_0		: 35
//PIN: ADDR_1		: 36
//PIN: ADDR_2		: 37
//PIN: ADDR_3		: 40
//PIN: ADDR_4		: 41
//PIN: ADDR_5		: 42
//PIN: ADDR_6		: 44
//PIN: ADDR_7		: 45
//PIN: ADDR_8		: 46
//PIN: ADDR_9		: 47
//PIN: ADDR_10		: 48
//PIN: ADDR_11		: 49
//PIN: ADDR_12		: 50
//PIN: ADDR_13		: 52
//PIN: ADDR_14		: 53
//PIN: ADDR_15		: 54
//PIN: ADDR_16		: 55
//PIN: ADDR_17		: 56
//PIN: ADDR_18		: 57
//PIN: ADDR_19		: 58
//PIN: ADDR_20		: 60
//PIN: ADDR_21		: 61
//PIN: ADDR_22		: 63
//PIN: ADDR_23		: 64
//PIN: ADDR_24		: 65
//PIN: ADDR_25		: 67
//PIN: ADDR_26		: 68
//PIN: ADDR_27		: 69
//PIN: ADDR_28		: 70
//PIN: ADDR_29		: 71
//PIN: ADDR_30		: 72
//PIN: ADDR_31		: 75
//PIN: FC_0		: 76
//PIN: FC_1		: 77
//PIN: FC_2		: 78
//PIN: nAS		: 87
//PIN: nDS		: 88
//PIN: nRST		: 89
//PIN: DRAM_CLK		: 90
//
//     === Outputs ===
//
//PIN: DSACK_0		: 1
//PIN: DSACK_1		: 2
//PIN: BERR		: 5
//PIN: CBACK		: 6
//PIN: STERM		: 7
//PIN: CI		: 8
//PIN: nFRAMSEL		: 9
//PIN: nFRAM_RD		: 10
//PIN: nFRAM_WR		: 12
//PIN: nFRAM_BE_0	: 13
//PIN: nFRAM_BE_1	: 14
//PIN: nFRAM_BE_2	: 16
//PIN: nFRAM_BE_3	: 17
//PIN: nEXPSEL		: 28
//PIN: nPSUCSEL		: 29
//PIN: nIACKSEL		: 79
//PIN: nINTCSEL		: 80
//PIN: nFPUSEL		: 81
//PIN: CPU_CLK		: 83
//PIN: CLK_6_25		: 84
//PIN: RESET		: 92
//PIN: nDRAMSEL_0	: 93
//PIN: nDRAMSEL_1	: 94
//PIN: nDRAMSEL_2	: 96
//PIN: nDRAMSEL_3	: 97
//PIN: nI2CSEL		: 98
//PIN: nISASEL		: 99
//PIN: nROMSEL		: 100
